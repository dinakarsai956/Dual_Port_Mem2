

package dual_port;
`include"packet.sv"
`include "transaction.sv"
//`include "interface.sv"
`include "generator.sv"
`include "driver.sv"
`include "driver_b.sv"
`include "monitor.sv"
`include "monitor_b.sv"
`include "reference.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include"test.sv"
endpackage : dual_port

